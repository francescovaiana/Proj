module norN1 #(parameter log_bit= 5) (in, out);
input [2**log_bit-1:0] in;
output out;

endmodule
